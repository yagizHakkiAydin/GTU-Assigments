module program_counter(
	output [31:0] pc_output,
	input [31:0] pc_input
);






endmodule