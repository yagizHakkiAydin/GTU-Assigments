module ONE_TO_32_EXTENDER(input inp , output [31:0] out);
	
	and a0(out[0],inp,inp);
	and a1(out[1],inp,inp);
	and a2(out[2],inp,inp);
	and a3(out[3],inp,inp);
	and a4(out[4],inp,inp);
	and a5(out[5],inp,inp);
	and a6(out[6],inp,inp);
	and a7(out[7],inp,inp);
	
	
	and a8(out[8],inp,inp);
	and a9(out[9],inp,inp);
	and a10(out[10],inp,inp);
	and a11(out[11],inp,inp);
	and a12(out[12],inp,inp);
	and a13(out[13],inp,inp);
	and a14(out[14],inp,inp);
	and a15(out[15],inp,inp);
	
	
	and a16(out[16],inp,inp);
	and a17(out[17],inp,inp);
	and a18(out[18],inp,inp);
	and a19(out[19],inp,inp);
	and a20(out[20],inp,inp);
	and a21(out[21],inp,inp);
	and a22(out[22],inp,inp);
	and a23(out[23],inp,inp);
	
	
	and a24(out[24],inp,inp);
	and a25(out[25],inp,inp);
	and a26(out[26],inp,inp);
	and a27(out[27],inp,inp);
	and a28(out[28],inp,inp);
	and a29(out[29],inp,inp);
	and a30(out[30],inp,inp);
	and a31(out[31],inp,inp);
	


endmodule




